/*******************************************************************
*
* Module: Memory.v
* Project: CSCE330_TermProject_MO
* Author: Mohamed Ashraf Taha - mohammedashraf@aucegypt.edu
          Omar Sherif Mahdy - omarmahdy122@aucegypt.edu
* Description: Combined memory that combines both instruction and data memories
*
* Change history: 04/23/20 - Combined data memory and instruction memory intoo one combined single memory that is byte addressable
*                          
*                 04/29/20 - Implemented the module as pipelined and combined memory
*                 05/03/20 - Decreased the capacity of the memory
*                 05/05/20 - fixed the bug of not loading from location of mem[0]
*                 05/06/20 - started testing sub cases of some functions to test the functionality of the memory and the full data_path
*                 05/09/20 
*                 05/10/20 
*                           - Full thorough testing of all the instructions
**********************************************************************/
`timescale 1ns / 1ps
module Memory
(input DmImSel,input clk, input MemRead, input MemWrite,
 input [2:0]Func3,
 input [31:0] addr, input [31:0] data_in,output reg [31:0] data_out);
 reg [7:0] mem [0:1023];
 wire [31:0] DataMemAddr;
 
assign DataMemAddr=  32'd1023-addr;

  always @(*) 
begin
    if (MemRead==1 && MemWrite==0 && DmImSel==0)
           begin
           case (Func3)
           3'b000: // LB
            data_out=mem[DataMemAddr];
            3'b001: // LH
             data_out={mem[DataMemAddr+1], mem[DataMemAddr]};
            3'b010: // LW
            begin
            if (addr==0)
            data_out= mem[DataMemAddr];
            else
             data_out={mem[DataMemAddr+3] ,mem[DataMemAddr+2],mem[DataMemAddr+1],mem[DataMemAddr]};
            end
            3'b100: //LBU
               data_out={{24{mem[DataMemAddr][7]}},mem[DataMemAddr]}; 
            3'b101: //LHU
            data_out = {{16{mem[DataMemAddr+1][7]}},mem[DataMemAddr+1],mem[DataMemAddr]};
           endcase
            end
    else if (MemWrite==1 && DmImSel==0)
           begin
           case (Func3[1:0])
           2'b00: //SB
             mem[DataMemAddr] = data_in[7:0];   
           2'b01:  //SH
               { mem[DataMemAddr+1],mem[DataMemAddr]} = data_in[15:0];   
           2'b10: // SW
                {mem[DataMemAddr+3] ,mem[DataMemAddr+2],mem[DataMemAddr+1],mem[DataMemAddr]} = data_in;   
           endcase
         
           end
           //INST MEM 
            else 
                      data_out= {mem[addr+3] ,mem[addr+2],mem[addr+1],mem[addr]};  
       end
//end


initial begin
{mem[1020],mem[1021],mem[1022],mem[1023]}=32'd10;// mem[0]
{mem[1016],mem[1017],mem[1018],mem[1019]}=32'd20;// mem[1]
{mem[1012],mem[1013],mem[1014],mem[1015]}=32'd30;    //mem[2]
{mem[1008],mem[1009],mem[1010],mem[1011]}=32'd40;    //mem[3]
{mem[1004],mem[1005],mem[1006],mem[1007]}=32'd50;    //mem[4]


 end
 
  initial begin
// OTHER INSTRUCTIONS TEST
               
//  {mem[3],mem[2],mem[1],mem[0]}=  32'b00000000110000110000001100010011; // addi  x6,x6,12               
//  {mem[7],mem[6],mem[5],mem[4]}=  32'b00000000000000000000011001100011; // Beq x0,x0,12 pc=4               
//  {mem[11],mem[10],mem[9],mem[8]}=  32'b00000000010100110000001010010011;//  addi x5,x6,5  8               
//  {mem[15],mem[14],mem[13],mem[12]}=  32'b00000000000100101100001000010011; // xori x4,x5,1 12               
//  {mem[19],mem[18],mem[17],mem[16]}=  32'b00000000000100100110000010010011; //ori x1, x4, 1 16               
//  {mem[23],mem[22],mem[21],mem[20]}=32'b000000000100_00000_010_00010_0000011 ; //lw x2, 4(x0)               
//  {mem[23],mem[22],mem[21],mem[20]}=32'b00000000011000000010011000100011 ; // sw x6, 16(x0)               
//  {mem[27],mem[26],mem[25],mem[24]}=32'b00000000000000000000000001110011;      //ecall          
//{mem[3],mem[2],mem[1],mem[0]}     =32'b0000000_00000_00000_000_00000_0110011;    // nop
//{mem[7],mem[6],mem[5],mem[4]}     =32'b00000000001000000000000010010011;    //addi x1,x0,2     // x1=2               
//{mem[11],mem[10],mem[9],mem[8]}   =32'b1111111_01100_00000_000_00010_0010011;    //addi x2,x0,-20   // x2= -20                                                     
//{mem[15],mem[14],mem[13],mem[12]} =32'b00000000011100000000000110010011;    //addi x3,x0,7     // x3=7//lw x3,0(x0)               
////{mem[15],mem[14],mem[13],mem[12]} =32'b00000000000000000010000110000011;     //lw x3,0(x0)               
//{mem[19],mem[18],mem[17],mem[16]} =32'b00000010000100011101011001100011;  // Bge x3,x1,44 , JUMP to ecall               
//////{mem[19],mem[18],mem[17],mem[16]} =32'b00000010000000000000011001100011;    // Beq x0,x0,44 , JUMP to ecall               
//{mem[23],mem[22],mem[21],mem[20]} =32'b11111111100000000000001000010011;    //addi x4,x0,-8    // x4= -8               
//{mem[27],mem[26],mem[25],mem[24]} =32'b01000000000100011000001010110011;    //sub x5, x3,x1    // x5= 5               
//{mem[31],mem[30],mem[29],mem[28]} =32'b01000000001100001000001100110011;    //sub x6, x1,x3    // x6= -5               
//{mem[35],mem[34],mem[33],mem[32]} =32'b01000000010000010000001110110011;    //sub x7, x2,x4 // x7=-12               
//{mem[39],mem[38],mem[37],mem[36]} =32'b01000000001100111000010000110011;    //sub x8, x7,x3 // x8= -19 	//FORWARDING CASE 1               
//{mem[43],mem[42],mem[41],mem[40]} =32'b01000000100000001000010010110011;    //sub x9, x1 ,x8 // x9=21  //FORWARDING CASE 2	               
//{mem[47],mem[46],mem[45],mem[44]} =32'b00000000000101001001010100010011;    //SLLI x10,x9,1 // x10=42  //FORWARDING CASE 3						               
//{mem[51],mem[50],mem[49],mem[48]} =32'b00000000000000000010010110000011;    //lw x11, 0(x0) // x11= 10               
//{mem[55],mem[54],mem[53],mem[52]} =32'b00000000000101011101011000010011;   	//SRLI x12,x11,1 // x12=5	//Load Use hazard CASE1S								               
//{mem[59],mem[58],mem[57],mem[56]} =32'b01000000000100100101011010010011;    //SRAI x13, x4, 1 //x13 = -4				                                
//{mem[63],mem[62],mem[61],mem[60]} = 32'b00000000000000000000000001110011;    //ecall                 
               
               
               
               
               
               
               
               
               
//{mem[3],mem[2],mem[1],mem[0]}          =32'b00000000000000000000000000110011         ;    //addi x0,x0,x0          
//{mem[7],mem[6],mem[5],mem[4]}          =32'b00000000001000000000000010010011         ;    //addi x1,x0,2           
//{mem[11],mem[10],mem[9],mem[8]}        =32'b11111110110000000000000100010011         ;    //addi x2,x0,-20         
//{mem[15],mem[14],mem[13],mem[12]}      =32'b00000000011100000000000110010011         ;    //addi x3,x0,7           
//{mem[19],mem[18],mem[17],mem[16]}      =32'b00000000011100000000000110010011         ;    //addi x4,x0,-8          
//{mem[23],mem[22],mem[21],mem[20]}      =32'b11111111100000000000001000010011         ;    //sub x5, x3,x1          
//{mem[27],mem[26],mem[25],mem[24]}      =32'b01000000000100011000001010110011         ;    //sub x6, x1,x3          
//{mem[31],mem[30],mem[29],mem[28]}      =32'b01000000001100001000001100110011         ;    //sub x7, x2,x4          
//{mem[35],mem[34],mem[33],mem[32]}      =32'b01000000010000010000001110110011         ;    //sub x8, x7,x3          
//{mem[39],mem[38],mem[37],mem[36]}      =32'b01000000001100111000010000110011         ;    //sub x9, x1 ,x8         
//{mem[43],mem[42],mem[41],mem[40]}      =32'b01000000100000001000010010110011         ;    //SLLI x10,x9,1          
//{mem[47],mem[46],mem[45],mem[44]}      =32'b00000000000101001001010100010011         ;    //lw x11, 0(x0)          
//{mem[51],mem[50],mem[49],mem[48]}      =32'b00000000000000000010010110000011         ;    //SRLI x12,x11,1         
//{mem[55],mem[54],mem[53],mem[52]}      =32'b00000000000101011101011000010011         ;    //SRAI x13,x4, 1         
//{mem[59],mem[58],mem[57],mem[56]}      =32'b01000000000100100101011010010000         ;    //andi x14,x5, 1         
//{mem[63],mem[62],mem[61],mem[60]}      =32'b00000000000100101111011100010011         ;    //andi x15,x5,-1         
//{mem[67],mem[66],mem[65],mem[64]}      =32'b11111111111100101111011110010011         ;    //ORI x16,x14,-2         
//{mem[71],mem[70],mem[69],mem[68]}      =32'b11111110011101110110100000010011         ;    //ORI x17,x14,25         
//{mem[75],mem[74],mem[73],mem[72]}      =32'b00000001100101110110100010010011         ;    //ORI x18,x2,-8          
//{mem[79],mem[78],mem[77],mem[76]}      =32'b00000000010000010110100100010011         ;    //Xor x19,x17,x1         
//{mem[83],mem[82],mem[81],mem[80]}      =32'b00000000000110001100100110110011         ;    //Xor x20,x2,x14         
//{mem[87],mem[86],mem[85],mem[84]}      =32'b00000000111000010100101000110011         ;    //Xor x21,x2,x7          
//{mem[91],mem[90],mem[89],mem[88]}      =32'b00000000011100010100101010110011         ;    //SLT x22,x1,x3          
//{mem[95],mem[94],mem[93],mem[92]}      =32'b00000000001100001010101100110011         ;    //SLT x23,x3,x1          
//{mem[99],mem[98],mem[97],mem[96]}      =32'b00000000000100011010101110110011         ;    //SLT x24,x4,x1          
//{mem[103],mem[102],mem[101],mem[100]}  =32'b00000000000100100010110000110011         ;    //SLT x25,x4,x6          
//{mem[107],mem[106],mem[105],mem[104]}  =32'b00000000011000100010110010110011         ;    //SLT x26,x6,x5          
//{mem[111],mem[110],mem[109],mem[108]}  =32'b00000000010100110010110100110011         ;    //SLT x27,x1,x4          
//{mem[115],mem[114],mem[113],mem[112]}  =32'b00000000010000001010110110110011         ;    //SLTu x28,x1,x3         
//{mem[119],mem[118],mem[117],mem[116]}  =32'b00000000001100001011111000110011         ;    //SLTu x29,x3,x1         
//{mem[123],mem[122],mem[121],mem[120]}  =32'b00000000000100011011111010110011         ;    //SLTu x30,x4,x1         
//{mem[127],mem[126],mem[125],mem[124]}  =32'b00000000000100100011111100110011         ;    //SLTu x31,x4,x6         
//{mem[131],mem[130],mem[129],mem[128]}  =32'b00000000011000100011111110110011         ;    //Xori x19,x17,2         
//{mem[131],mem[130],mem[129],mem[128]}  =32'b00000000000000000000000110000011         ;    //Xori x20,x2,1          
//{mem[135],mem[134],mem[133],mem[132]}  =32'b01111111011000011000001000010011         ;    //Xori x21,x2,-1         
//{mem[139],mem[138],mem[137],mem[136]}  =32'b00000000010000000010110000100011         ;    //SLTu x1,x6,x5          
//{mem[143],mem[142],mem[141],mem[140]}  =32'b00000000010000000001111000100011         ;    //SLTu x2,x1,x4 
////{mem[147],mem[146],mem[145],mem[144]} =32'b00000000000000000000000001110011 ;           //ecall     
//{mem[147],mem[146],mem[145],mem[144]}  =32'b00000000000000000000000110000011         ;    // #lb x3,0(x0)   
//{mem[151],mem[150],mem[149],mem[148]}  =32'b01111111011000011000001000010011         ;    // addi x4,x3,2038
//{mem[155],mem[154],mem[153],mem[152]}  =32'b00000000010000000010110000100011         ;    // #sw x4,24(x0)  
//{mem[159],mem[158],mem[157],mem[156]}  =32'b00000000010000000001111000100011         ;    // #sh x4,28(x0)  
//{mem[163],mem[162],mem[161],mem[160]}  =32'b00001000000100000000001010010011         ;    // addi x5,x0,129 
//{mem[167],mem[166],mem[165],mem[164]}  =32'b00000010010100000001000000100011         ;    // #sh x5,32(x0)	   
//{mem[171],mem[170],mem[169],mem[168]}  =32'b00000010010100000000001000100011         ;    // #sb x5,36(x0)	     
//{mem[175],mem[174],mem[173],mem[172]}  =32'b10000000000000000000001100010011         ;    // addi x6,x0,-327
//{mem[179],mem[178],mem[177],mem[176]}  =32'b11110111111100000000001110010011         ;    // addi x7,x0,-129
//{mem[183],mem[182],mem[181],mem[180]}  =32'b00000010011000000010010000100011         ;    // #sw x6,40(x0)  
//{mem[187],mem[186],mem[185],mem[184]}  =32'b00000010011000000001011000100011         ;    // #sh x6,44(x0)  
//{mem[191],mem[190],mem[189],mem[188]}  =32'b00000010011100000001100000100011         ;    // #sh x7,48(x0)	     
//{mem[195],mem[194],mem[193],mem[192]}  =32'b00000010011100000000101000100011         ;    // #sb x7,52(x0)	     
//{mem[199],mem[198],mem[197],mem[196]}  =32'b00000001100000000001010000000011         ;    // #lh x8,24(x0)	     
//{mem[203],mem[202],mem[201],mem[200]}  =32'b00000001100000000010010010000011         ;    // #lw x9,24(x0)  
//{mem[207],mem[206],mem[205],mem[204]}  =32'b00000010000000000001010100000011         ;    // #lh x10,32(x0)	   
//{mem[211],mem[210],mem[209],mem[208]}  =32'b00000010000000000000010110000011         ;    // #lb x11,32(x0) 
//{mem[215],mem[214],mem[213],mem[212]}  =32'b00000010100000000001011000000011         ;    // #lh x12,40(x0)	   
//{mem[219],mem[218],mem[217],mem[216]}  =32'b00000010100000000101011010000011         ;    // #lhu x13,40(x0)
//{mem[223],mem[222],mem[221],mem[220]}  =32'b00000011000000000000011100000011         ;    // #lb x14,48(x0)	            
//{mem[227],mem[226],mem[225],mem[224]}  =32'b00000011000000000100011110000011         ;    // #lbu x15,48(x0)
//{mem[231],mem[230],mem[229],mem[228]}  =32'b00000000001000100110100000110111         ;    // lui x16, 550   
//{mem[235],mem[234],mem[233],mem[232]}  =32'b00000000010100000000100010010011         ;    // addi x17,x0,5  
//{mem[239],mem[238],mem[237],mem[236]}  =32'b00000000010100000000100100010011         ;    // addi x18, x0,5 
//{mem[243],mem[242],mem[241],mem[240]}  =32'b00000000000000000000000001110011          ;   //ecall  
     
                                                                                                                      
//BRANCH TEST




//{mem[3],mem[2],mem[1],mem[0]}          =32'b00000000000000000000000000010011;  //addi x0,x0,x0          
//{mem[7],mem[6],mem[5],mem[4]}          =32'b00000000000000000010000010000011;  //lw x1,0(x0)          
//{mem[11],mem[10],mem[9],mem[8]}        =32'b00000000001000001101110001100011;  //addi x2,x0,3         
//{mem[15],mem[14],mem[13],mem[12]}      =32'b00000000000000000000000000010011;  //bge x1,x2,20                 
//{mem[19],mem[18],mem[17],mem[16]}      =32'b00000000000000000000000000010011;  //nop	         
//{mem[23],mem[22],mem[21],mem[20]}      =32'b00000000000000000000000000010011;  //nop	        
//{mem[27],mem[26],mem[25],mem[24]}      =32'b00000000000000000000000000010011;  //nop	        
//{mem[31],mem[30],mem[29],mem[28]}      =32'b00000000000100010000000110110011;  //add x3,x2,x1
//{mem[35],mem[34],mem[33],mem[32]}      =32'b00000000001100001101110001100011;  //bge x1,x3,20 
//{mem[39],mem[38],mem[37],mem[36]}      =32'b00000010001100001100100001100011;  //blt x1,x3,44
//{mem[43],mem[42],mem[41],mem[40]}      =32'b00000000000000000000000000010011;   //nop       
//{mem[47],mem[46],mem[45],mem[44]}      =32'b00000000000000000000000000010011;   //nop       
//{mem[51],mem[50],mem[49],mem[48]}      =32'b00000000000000000000000000010011;   //nop       
//{mem[55],mem[54],mem[53],mem[52]}      =32'b00000000000000000000000000010011;   //nop       
//{mem[59],mem[58],mem[57],mem[56]}      =32'b00000000000000000000000000010011;   //nop       
//{mem[63],mem[62],mem[61],mem[60]}      =32'b00000000000000000000000000010011;   //nop       
//{mem[67],mem[66],mem[65],mem[64]}      =32'b00000000000000000000000000010011;   //nop       
//{mem[71],mem[70],mem[69],mem[68]}      =32'b00000000000000000000000000010011;   //nop       
//{mem[75],mem[74],mem[73],mem[72]}      =32'b00000000000000000000000000010011;   //nop       
//{mem[79],mem[78],mem[77],mem[76]}      =32'b00000000000000000000000000010011;   //nop       
//{mem[83],mem[82],mem[81],mem[80]}      =32'b00000000101000000000000100010011;   //addi x2,x0,10      
//{mem[87],mem[86],mem[85],mem[84]}      =32'b00000000001100010001100101100011;   //blt x3,x2, 40        
//{mem[91],mem[90],mem[89],mem[88]}      =32'b00000010001000011100010001100011;   //beq x2,x3, 16 
//{mem[95],mem[94],mem[93],mem[92]}      =32'b00000000001100010000100001100011;     //nop
//{mem[99],mem[98],mem[97],mem[96]}      =32'b00000000000000000000000000010011;     //nop
//{mem[103],mem[102],mem[101],mem[100]}  =32'b00000000000000000000000000010011;     //nop
//{mem[107],mem[106],mem[105],mem[104]}  =32'b00000000000000000000000000010011;     //nop
//{mem[111],mem[110],mem[109],mem[108]}  =32'b00000010010000010000001001100011;    //addi x4,x0,10
//{mem[115],mem[114],mem[113],mem[112]}  =32'b00000000010000010001110001100011;   //beq x2,x4, 32
//{mem[119],mem[118],mem[117],mem[116]}  =32'b00000000010000010001101001100011;   //bne x2,x4,20
//{mem[123],mem[122],mem[121],mem[120]}  =32'b00000000000000000000000000010011;    //nop
//{mem[127],mem[126],mem[125],mem[124]}  =32'b00000000000000000000000000010011;    //nop
//{mem[131],mem[130],mem[129],mem[128]}  =32'b00000000000000000000000000010011;    //nop
//{mem[135],mem[134],mem[133],mem[132]}  =32'b00000000000000000000000000010011;    //nop
//{mem[139],mem[138],mem[137],mem[136]}  =32'b00000000001100010001100101100011;   //bne x2,x13,0 NT	    
//{mem[143],mem[142],mem[141],mem[140]}=32'b00000000000000000000000001110011;   //ecall 

                                          
                                                                                        


 {mem[3],mem[2],mem[1],mem[0]}    =32'b00000000000000000000000000010011;  //addi x0,x0,x0
 {mem[7],mem[6],mem[5],mem[4]}    = 32'b00000000000000000010000010000011 ;//lw x1,0(x0)               x1=10
 {mem[11],mem[10],mem[9],mem[8]}  = 32'b00000000001100000000000100010011 ;//addi x2,x0,3              x2=3
 {mem[15],mem[14],mem[13],mem[12]}= 32'b00000010000100010000000110110011 ;// mul x3,x2,x1             x3=30
 {mem[19],mem[18],mem[17],mem[16]}= 32'b00000010000100010001001000110011 ;// mulh x4,x2,x1            x4= ???
 {mem[23],mem[22],mem[21],mem[20]}= 32'b00000010000100010010001010110011 ;// mulhsu x5,x2,x1          x5=??
 {mem[27],mem[26],mem[25],mem[24]}= 32'b00000010000100010011001100110011 ;// mulhu x6,x2,x1           x6=?    
 {mem[31],mem[30],mem[29],mem[28]}= 32'b00000010000100011100001110110011 ;// DIV x7,x3,x1             x7 = 3
 {mem[35],mem[34],mem[33],mem[32]}= 32'b11111111010000000000010000010011 ;// addi x8,x0,-12           x8=-12
 {mem[39],mem[38],mem[37],mem[36]}= 32'b00000010000101000101010010110011 ;// DIVU x9, x8, x1          x9 =????
 {mem[43],mem[42],mem[41],mem[40]}= 32'b00000010001100001110010100110011 ;// rem x10, x1,x3           x10=1
 {mem[47],mem[46],mem[45],mem[44]}= 32'b00000010001101000111010110110011 ;// remu x11,x8,x3           x11=??
 {mem[51],mem[50],mem[49],mem[48]}  =32'b00000000000000000000000001110011;   //ecall 
 
 
 
 
 
 
 
  end                                              
                                                   
 
endmodule                                                                   





 
 

   
   
   

 
 
   
   
   
 
  
 
  
 
  
 



                    
                    
                    
                    
                    
                    
                    
                    
                    
                    
                    
                    
                    
                    
                    
                    
                    
                    































